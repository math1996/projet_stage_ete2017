----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:34:40 07/18/2017 
-- Design Name: 
-- Module Name:    LUT_256_gain - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LUT_256_gain is
    Port ( adresse : in  STD_LOGIC_VECTOR (7 downto 0);
           valeur : out  STD_LOGIC_VECTOR (31 downto 0));
end LUT_256_gain;

architecture Behavioral of LUT_256_gain is

begin

process(adresse)
begin
	case adresse is
		when "00000000" => valeur <="01111111111111111111111111111111";
		when "00000001" => valeur <="00000001000000110110101110111010";
		when "00000010" => valeur <="00000000100000011011010111011101";
		when "00000011" => valeur <="00000000010101100111100100111110";
		when "00000100" => valeur <="00000000010000001101101011101111";
		when "00000101" => valeur <="00000000001100111110001001011000";
		when "00000110" => valeur <="00000000001010110011110010011111";
		when "00000111" => valeur <="00000000001001010000111101100100";
		when "00001000" => valeur <="00000000001000000110110101110111";
		when "00001001" => valeur <="00000000000111001101001100010101";
		when "00001010" => valeur <="00000000000110011111000100101100";
		when "00001011" => valeur <="00000000000101111001010101101110";
		when "00001100" => valeur <="00000000000101011001111001010000";
		when "00001101" => valeur <="00000000000100111111010010011000";
		when "00001110" => valeur <="00000000000100101000011110110010";
		when "00001111" => valeur <="00000000000100010100101101110011";
		when "00010000" => valeur <="00000000000100000011011010111100";
		when "00010001" => valeur <="00000000000011110100001010010010";
		when "00010010" => valeur <="00000000000011100110100110001010";
		when "00010011" => valeur <="00000000000011011010011101011011";
		when "00010100" => valeur <="00000000000011001111100010010110";
		when "00010101" => valeur <="00000000000011000101101001110111";
		when "00010110" => valeur <="00000000000010111100101010110111";
		when "00010111" => valeur <="00000000000010110100011101110111";
		when "00011000" => valeur <="00000000000010101100111100101000";
		when "00011001" => valeur <="00000000000010100110000001111000";
		when "00011010" => valeur <="00000000000010011111101001001100";
		when "00011011" => valeur <="00000000000010011001101110110010";
		when "00011100" => valeur <="00000000000010010100001111011001";
		when "00011101" => valeur <="00000000000010001111001000001111";
		when "00011110" => valeur <="00000000000010001010010110111001";
		when "00011111" => valeur <="00000000000010000101111001010000";
		when "00100000" => valeur <="00000000000010000001101101011110";
		when "00100001" => valeur <="00000000000001111101110001111010";
		when "00100010" => valeur <="00000000000001111010000101001001";
		when "00100011" => valeur <="00000000000001110110100101111010";
		when "00100100" => valeur <="00000000000001110011010011000101";
		when "00100101" => valeur <="00000000000001110000001011101001";
		when "00100110" => valeur <="00000000000001101101001110101101";
		when "00100111" => valeur <="00000000000001101010011011011101";
		when "00101000" => valeur <="00000000000001100111110001001011";
		when "00101001" => valeur <="00000000000001100101001111001100";
		when "00101010" => valeur <="00000000000001100010110100111011";
		when "00101011" => valeur <="00000000000001100000100001110101";
		when "00101100" => valeur <="00000000000001011110010101011100";
		when "00101101" => valeur <="00000000000001011100001111010001";
		when "00101110" => valeur <="00000000000001011010001110111100";
		when "00101111" => valeur <="00000000000001011000010100000100";
		when "00110000" => valeur <="00000000000001010110011110010100";
		when "00110001" => valeur <="00000000000001010100101101010111";
		when "00110010" => valeur <="00000000000001010011000000111100";
		when "00110011" => valeur <="00000000000001010001011000110001";
		when "00110100" => valeur <="00000000000001001111110100100110";
		when "00110101" => valeur <="00000000000001001110010100001101";
		when "00110110" => valeur <="00000000000001001100110111011001";
		when "00110111" => valeur <="00000000000001001011011101111100";
		when "00111000" => valeur <="00000000000001001010000111101100";
		when "00111001" => valeur <="00000000000001001000110100011110";
		when "00111010" => valeur <="00000000000001000111100100001000";
		when "00111011" => valeur <="00000000000001000110010110011111";
		when "00111100" => valeur <="00000000000001000101001011011101";
		when "00111101" => valeur <="00000000000001000100000010111000";
		when "00111110" => valeur <="00000000000001000010111100101000";
		when "00111111" => valeur <="00000000000001000001111000101000";
		when "01000000" => valeur <="00000000000001000000110110101111";
		when "01000001" => valeur <="00000000000000111111110110111000";
		when "01000010" => valeur <="00000000000000111110111000111101";
		when "01000011" => valeur <="00000000000000111101111100111000";
		when "01000100" => valeur <="00000000000000111101000010100101";
		when "01000101" => valeur <="00000000000000111100001001111101";
		when "01000110" => valeur <="00000000000000111011010010111101";
		when "01000111" => valeur <="00000000000000111010011101100000";
		when "01001000" => valeur <="00000000000000111001101001100011";
		when "01001001" => valeur <="00000000000000111000110111000000";
		when "01001010" => valeur <="00000000000000111000000101110101";
		when "01001011" => valeur <="00000000000000110111010101111101";
		when "01001100" => valeur <="00000000000000110110100111010111";
		when "01001101" => valeur <="00000000000000110101111001111101";
		when "01001110" => valeur <="00000000000000110101001101101111";
		when "01001111" => valeur <="00000000000000110100100010101000";
		when "01010000" => valeur <="00000000000000110011111000100110";
		when "01010001" => valeur <="00000000000000110011001111100110";
		when "01010010" => valeur <="00000000000000110010100111100110";
		when "01010011" => valeur <="00000000000000110010000000100100";
		when "01010100" => valeur <="00000000000000110001011010011110";
		when "01010101" => valeur <="00000000000000110000110101010000";
		when "01010110" => valeur <="00000000000000110000010000111011";
		when "01010111" => valeur <="00000000000000101111101101011010";
		when "01011000" => valeur <="00000000000000101111001010101110";
		when "01011001" => valeur <="00000000000000101110101000110011";
		when "01011010" => valeur <="00000000000000101110000111101000";
		when "01011011" => valeur <="00000000000000101101100111001101";
		when "01011100" => valeur <="00000000000000101101000111011110";
		when "01011101" => valeur <="00000000000000101100101000011011";
		when "01011110" => valeur <="00000000000000101100001010000010";
		when "01011111" => valeur <="00000000000000101011101100010010";
		when "01100000" => valeur <="00000000000000101011001111001010";
		when "01100001" => valeur <="00000000000000101010110010101000";
		when "01100010" => valeur <="00000000000000101010010110101100";
		when "01100011" => valeur <="00000000000000101001111011010011";
		when "01100100" => valeur <="00000000000000101001100000011110";
		when "01100101" => valeur <="00000000000000101001000110001011";
		when "01100110" => valeur <="00000000000000101000101100011000";
		when "01100111" => valeur <="00000000000000101000010011000110";
		when "01101000" => valeur <="00000000000000100111111010010011";
		when "01101001" => valeur <="00000000000000100111100001111110";
		when "01101010" => valeur <="00000000000000100111001010000111";
		when "01101011" => valeur <="00000000000000100110110010101100";
		when "01101100" => valeur <="00000000000000100110011011101100";
		when "01101101" => valeur <="00000000000000100110000101001000";
		when "01101110" => valeur <="00000000000000100101101110111110";
		when "01101111" => valeur <="00000000000000100101011001001110";
		when "01110000" => valeur <="00000000000000100101000011110110";
		when "01110001" => valeur <="00000000000000100100101110110111";
		when "01110010" => valeur <="00000000000000100100011010001111";
		when "01110011" => valeur <="00000000000000100100000101111110";
		when "01110100" => valeur <="00000000000000100011110010000100";
		when "01110101" => valeur <="00000000000000100011011110011111";
		when "01110110" => valeur <="00000000000000100011001011010000";
		when "01110111" => valeur <="00000000000000100010111000010101";
		when "01111000" => valeur <="00000000000000100010100101101110";
		when "01111001" => valeur <="00000000000000100010010011011011";
		when "01111010" => valeur <="00000000000000100010000001011100";
		when "01111011" => valeur <="00000000000000100001101111101111";
		when "01111100" => valeur <="00000000000000100001011110010100";
		when "01111101" => valeur <="00000000000000100001001101001011";
		when "01111110" => valeur <="00000000000000100000111100010100";
		when "01111111" => valeur <="00000000000000100000101011101101";
		when "10000000" => valeur <="00000000000000100000011011010111";
		when "10000001" => valeur <="00000000000000100000001011010010";
		when "10000010" => valeur <="00000000000000011111111011011100";
		when "10000011" => valeur <="00000000000000011111101011110110";
		when "10000100" => valeur <="00000000000000011111011100011111";
		when "10000101" => valeur <="00000000000000011111001101010110";
		when "10000110" => valeur <="00000000000000011110111110011100";
		when "10000111" => valeur <="00000000000000011110101111110000";
		when "10001000" => valeur <="00000000000000011110100001010010";
		when "10001001" => valeur <="00000000000000011110010011000010";
		when "10001010" => valeur <="00000000000000011110000100111111";
		when "10001011" => valeur <="00000000000000011101110111001000";
		when "10001100" => valeur <="00000000000000011101101001011111";
		when "10001101" => valeur <="00000000000000011101011100000001";
		when "10001110" => valeur <="00000000000000011101001110110000";
		when "10001111" => valeur <="00000000000000011101000001101011";
		when "10010000" => valeur <="00000000000000011100110100110001";
		when "10010001" => valeur <="00000000000000011100101000000011";
		when "10010010" => valeur <="00000000000000011100011011100000";
		when "10010011" => valeur <="00000000000000011100001111001000";
		when "10010100" => valeur <="00000000000000011100000010111010";
		when "10010101" => valeur <="00000000000000011011110110110111";
		when "10010110" => valeur <="00000000000000011011101010111111";
		when "10010111" => valeur <="00000000000000011011011111010000";
		when "10011000" => valeur <="00000000000000011011010011101011";
		when "10011001" => valeur <="00000000000000011011001000010000";
		when "10011010" => valeur <="00000000000000011010111100111111";
		when "10011011" => valeur <="00000000000000011010110001110110";
		when "10011100" => valeur <="00000000000000011010100110110111";
		when "10011101" => valeur <="00000000000000011010011100000001";
		when "10011110" => valeur <="00000000000000011010010001010100";
		when "10011111" => valeur <="00000000000000011010000110101111";
		when "10100000" => valeur <="00000000000000011001111100010011";
		when "10100001" => valeur <="00000000000000011001110001111111";
		when "10100010" => valeur <="00000000000000011001100111110011";
		when "10100011" => valeur <="00000000000000011001011101101111";
		when "10100100" => valeur <="00000000000000011001010011110011";
		when "10100101" => valeur <="00000000000000011001001001111111";
		when "10100110" => valeur <="00000000000000011001000000010010";
		when "10100111" => valeur <="00000000000000011000110110101101";
		when "10101000" => valeur <="00000000000000011000101101001111";
		when "10101001" => valeur <="00000000000000011000100011111000";
		when "10101010" => valeur <="00000000000000011000011010101000";
		when "10101011" => valeur <="00000000000000011000010001011111";
		when "10101100" => valeur <="00000000000000011000001000011101";
		when "10101101" => valeur <="00000000000000010111111111100010";
		when "10101110" => valeur <="00000000000000010111110110101101";
		when "10101111" => valeur <="00000000000000010111101101111111";
		when "10110000" => valeur <="00000000000000010111100101010111";
		when "10110001" => valeur <="00000000000000010111011100110101";
		when "10110010" => valeur <="00000000000000010111010100011001";
		when "10110011" => valeur <="00000000000000010111001100000100";
		when "10110100" => valeur <="00000000000000010111000011110100";
		when "10110101" => valeur <="00000000000000010110111011101010";
		when "10110110" => valeur <="00000000000000010110110011100110";
		when "10110111" => valeur <="00000000000000010110101011101000";
		when "10111000" => valeur <="00000000000000010110100011101111";
		when "10111001" => valeur <="00000000000000010110011011111011";
		when "10111010" => valeur <="00000000000000010110010100001101";
		when "10111011" => valeur <="00000000000000010110001100100101";
		when "10111100" => valeur <="00000000000000010110000101000001";
		when "10111101" => valeur <="00000000000000010101111101100011";
		when "10111110" => valeur <="00000000000000010101110110001001";
		when "10111111" => valeur <="00000000000000010101101110110101";
		when "11000000" => valeur <="00000000000000010101100111100101";
		when "11000001" => valeur <="00000000000000010101100000011010";
		when "11000010" => valeur <="00000000000000010101011001010100";
		when "11000011" => valeur <="00000000000000010101010010010011";
		when "11000100" => valeur <="00000000000000010101001011010110";
		when "11000101" => valeur <="00000000000000010101000100011110";
		when "11000110" => valeur <="00000000000000010100111101101010";
		when "11000111" => valeur <="00000000000000010100110110111010";
		when "11001000" => valeur <="00000000000000010100110000001111";
		when "11001001" => valeur <="00000000000000010100101001101000";
		when "11001010" => valeur <="00000000000000010100100011000101";
		when "11001011" => valeur <="00000000000000010100011100100111";
		when "11001100" => valeur <="00000000000000010100010110001100";
		when "11001101" => valeur <="00000000000000010100001111110110";
		when "11001110" => valeur <="00000000000000010100001001100011";
		when "11001111" => valeur <="00000000000000010100000011010100";
		when "11010000" => valeur <="00000000000000010011111101001010";
		when "11010001" => valeur <="00000000000000010011110111000010";
		when "11010010" => valeur <="00000000000000010011110000111111";
		when "11010011" => valeur <="00000000000000010011101010111111";
		when "11010100" => valeur <="00000000000000010011100101000011";
		when "11010101" => valeur <="00000000000000010011011111001011";
		when "11010110" => valeur <="00000000000000010011011001010110";
		when "11010111" => valeur <="00000000000000010011010011100100";
		when "11011000" => valeur <="00000000000000010011001101110110";
		when "11011001" => valeur <="00000000000000010011001000001011";
		when "11011010" => valeur <="00000000000000010011000010100100";
		when "11011011" => valeur <="00000000000000010010111101000000";
		when "11011100" => valeur <="00000000000000010010110111011111";
		when "11011101" => valeur <="00000000000000010010110010000001";
		when "11011110" => valeur <="00000000000000010010101100100111";
		when "11011111" => valeur <="00000000000000010010100111001111";
		when "11100000" => valeur <="00000000000000010010100001111011";
		when "11100001" => valeur <="00000000000000010010011100101010";
		when "11100010" => valeur <="00000000000000010010010111011011";
		when "11100011" => valeur <="00000000000000010010010010010000";
		when "11100100" => valeur <="00000000000000010010001101001000";
		when "11100101" => valeur <="00000000000000010010001000000010";
		when "11100110" => valeur <="00000000000000010010000010111111";
		when "11100111" => valeur <="00000000000000010001111101111111";
		when "11101000" => valeur <="00000000000000010001111001000010";
		when "11101001" => valeur <="00000000000000010001110100000111";
		when "11101010" => valeur <="00000000000000010001101111010000";
		when "11101011" => valeur <="00000000000000010001101010011010";
		when "11101100" => valeur <="00000000000000010001100101101000";
		when "11101101" => valeur <="00000000000000010001100000111000";
		when "11101110" => valeur <="00000000000000010001011100001010";
		when "11101111" => valeur <="00000000000000010001010111100000";
		when "11110000" => valeur <="00000000000000010001010010110111";
		when "11110001" => valeur <="00000000000000010001001110010001";
		when "11110010" => valeur <="00000000000000010001001001101110";
		when "11110011" => valeur <="00000000000000010001000101001101";
		when "11110100" => valeur <="00000000000000010001000000101110";
		when "11110101" => valeur <="00000000000000010000111100010001";
		when "11110110" => valeur <="00000000000000010000110111110111";
		when "11110111" => valeur <="00000000000000010000110011100000";
		when "11111000" => valeur <="00000000000000010000101111001010";
		when "11111001" => valeur <="00000000000000010000101010110111";
		when "11111010" => valeur <="00000000000000010000100110100110";
		when "11111011" => valeur <="00000000000000010000100010010111";
		when "11111100" => valeur <="00000000000000010000011110001010";
		when "11111101" => valeur <="00000000000000010000011001111111";
		when "11111110" => valeur <="00000000000000010000010101110111";
		when "11111111" => valeur <="00000000000000010000010001110000";
		when others => valeur <= (others => '0');
	end case;
end process;

end Behavioral;

