----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    09:51:54 05/30/2017 
-- Design Name: 
-- Module Name:    LUT_1024_sin - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity LUT_1024_sin is
    Port ( adresse : in  STD_LOGIC_VECTOR (9 downto 0);
           valeur : out  STD_LOGIC_VECTOR (15 downto 0));
end LUT_1024_sin;

architecture Behavioral of LUT_1024_sin is

begin

process(adresse)
begin
	case adresse is 
		when "0000000000" => valeur <= X"0000";
		when "0000000001" => valeur <= X"0016";
		when "0000000010" => valeur <= X"002C";
		when "0000000011" => valeur <= X"0042";
		when "0000000100" => valeur <= X"0057";
		when "0000000101" => valeur <= X"006D";
		when "0000000110" => valeur <= X"0083";
		when "0000000111" => valeur <= X"0099";
		when "0000001000" => valeur <= X"00AF";
		when "0000001001" => valeur <= X"00C5";
		when "0000001010" => valeur <= X"00DB";
		when "0000001011" => valeur <= X"00F0";
		when "0000001100" => valeur <= X"0106";
		when "0000001101" => valeur <= X"011C";
		when "0000001110" => valeur <= X"0132";
		when "0000001111" => valeur <= X"0148";
		when "0000010000" => valeur <= X"015E";
		when "0000010001" => valeur <= X"0174";
		when "0000010010" => valeur <= X"0189";
		when "0000010011" => valeur <= X"019F";
		when "0000010100" => valeur <= X"01B5";
		when "0000010101" => valeur <= X"01CB";
		when "0000010110" => valeur <= X"01E1";
		when "0000010111" => valeur <= X"01F6";
		when "0000011000" => valeur <= X"020C";
		when "0000011001" => valeur <= X"0222";
		when "0000011010" => valeur <= X"0238";
		when "0000011011" => valeur <= X"024E";
		when "0000011100" => valeur <= X"0263";
		when "0000011101" => valeur <= X"0279";
		when "0000011110" => valeur <= X"028F";
		when "0000011111" => valeur <= X"02A5";
		when "0000100000" => valeur <= X"02BB";
		when "0000100001" => valeur <= X"02D0";
		when "0000100010" => valeur <= X"02E6";
		when "0000100011" => valeur <= X"02FC";
		when "0000100100" => valeur <= X"0311";
		when "0000100101" => valeur <= X"0327";
		when "0000100110" => valeur <= X"033D";
		when "0000100111" => valeur <= X"0353";
		when "0000101000" => valeur <= X"0368";
		when "0000101001" => valeur <= X"037E";
		when "0000101010" => valeur <= X"0394";
		when "0000101011" => valeur <= X"03A9";
		when "0000101100" => valeur <= X"03BF";
		when "0000101101" => valeur <= X"03D5";
		when "0000101110" => valeur <= X"03EA";
		when "0000101111" => valeur <= X"0400";
		when "0000110000" => valeur <= X"0416";
		when "0000110001" => valeur <= X"042B";
		when "0000110010" => valeur <= X"0441";
		when "0000110011" => valeur <= X"0457";
		when "0000110100" => valeur <= X"046C";
		when "0000110101" => valeur <= X"0482";
		when "0000110110" => valeur <= X"0497";
		when "0000110111" => valeur <= X"04AD";
		when "0000111000" => valeur <= X"04C2";
		when "0000111001" => valeur <= X"04D8";
		when "0000111010" => valeur <= X"04ED";
		when "0000111011" => valeur <= X"0503";
		when "0000111100" => valeur <= X"0518";
		when "0000111101" => valeur <= X"052E";
		when "0000111110" => valeur <= X"0543";
		when "0000111111" => valeur <= X"0559";
		when "0001000000" => valeur <= X"056E";
		when "0001000001" => valeur <= X"0584";
		when "0001000010" => valeur <= X"0599";
		when "0001000011" => valeur <= X"05AF";
		when "0001000100" => valeur <= X"05C4";
		when "0001000101" => valeur <= X"05D9";
		when "0001000110" => valeur <= X"05EF";
		when "0001000111" => valeur <= X"0604";
		when "0001001000" => valeur <= X"0619";
		when "0001001001" => valeur <= X"062F";
		when "0001001010" => valeur <= X"0644";
		when "0001001011" => valeur <= X"0659";
		when "0001001100" => valeur <= X"066F";
		when "0001001101" => valeur <= X"0684";
		when "0001001110" => valeur <= X"0699";
		when "0001001111" => valeur <= X"06AE";
		when "0001010000" => valeur <= X"06C4";
		when "0001010001" => valeur <= X"06D9";
		when "0001010010" => valeur <= X"06EE";
		when "0001010011" => valeur <= X"0703";
		when "0001010100" => valeur <= X"0718";
		when "0001010101" => valeur <= X"072D";
		when "0001010110" => valeur <= X"0743";
		when "0001010111" => valeur <= X"0758";
		when "0001011000" => valeur <= X"076D";
		when "0001011001" => valeur <= X"0782";
		when "0001011010" => valeur <= X"0797";
		when "0001011011" => valeur <= X"07AC";
		when "0001011100" => valeur <= X"07C1";
		when "0001011101" => valeur <= X"07D6";
		when "0001011110" => valeur <= X"07EB";
		when "0001011111" => valeur <= X"0800";
		when "0001100000" => valeur <= X"0815";
		when "0001100001" => valeur <= X"082A";
		when "0001100010" => valeur <= X"083E";
		when "0001100011" => valeur <= X"0853";
		when "0001100100" => valeur <= X"0868";
		when "0001100101" => valeur <= X"087D";
		when "0001100110" => valeur <= X"0892";
		when "0001100111" => valeur <= X"08A7";
		when "0001101000" => valeur <= X"08BB";
		when "0001101001" => valeur <= X"08D0";
		when "0001101010" => valeur <= X"08E5";
		when "0001101011" => valeur <= X"08FA";
		when "0001101100" => valeur <= X"090E";
		when "0001101101" => valeur <= X"0923";
		when "0001101110" => valeur <= X"0938";
		when "0001101111" => valeur <= X"094C";
		when "0001110000" => valeur <= X"0961";
		when "0001110001" => valeur <= X"0975";
		when "0001110010" => valeur <= X"098A";
		when "0001110011" => valeur <= X"099E";
		when "0001110100" => valeur <= X"09B3";
		when "0001110101" => valeur <= X"09C7";
		when "0001110110" => valeur <= X"09DC";
		when "0001110111" => valeur <= X"09F0";
		when "0001111000" => valeur <= X"0A05";
		when "0001111001" => valeur <= X"0A19";
		when "0001111010" => valeur <= X"0A2D";
		when "0001111011" => valeur <= X"0A42";
		when "0001111100" => valeur <= X"0A56";
		when "0001111101" => valeur <= X"0A6A";
		when "0001111110" => valeur <= X"0A7F";
		when "0001111111" => valeur <= X"0A93";
		when "0010000000" => valeur <= X"0AA7";
		when "0010000001" => valeur <= X"0ABB";
		when "0010000010" => valeur <= X"0ACF";
		when "0010000011" => valeur <= X"0AE4";
		when "0010000100" => valeur <= X"0AF8";
		when "0010000101" => valeur <= X"0B0C";
		when "0010000110" => valeur <= X"0B20";
		when "0010000111" => valeur <= X"0B34";
		when "0010001000" => valeur <= X"0B48";
		when "0010001001" => valeur <= X"0B5C";
		when "0010001010" => valeur <= X"0B70";
		when "0010001011" => valeur <= X"0B84";
		when "0010001100" => valeur <= X"0B98";
		when "0010001101" => valeur <= X"0BAB";
		when "0010001110" => valeur <= X"0BBF";
		when "0010001111" => valeur <= X"0BD3";
		when "0010010000" => valeur <= X"0BE7";
		when "0010010001" => valeur <= X"0BFB";
		when "0010010010" => valeur <= X"0C0E";
		when "0010010011" => valeur <= X"0C22";
		when "0010010100" => valeur <= X"0C36";
		when "0010010101" => valeur <= X"0C49";
		when "0010010110" => valeur <= X"0C5D";
		when "0010010111" => valeur <= X"0C70";
		when "0010011000" => valeur <= X"0C84";
		when "0010011001" => valeur <= X"0C98";
		when "0010011010" => valeur <= X"0CAB";
		when "0010011011" => valeur <= X"0CBE";
		when "0010011100" => valeur <= X"0CD2";
		when "0010011101" => valeur <= X"0CE5";
		when "0010011110" => valeur <= X"0CF9";
		when "0010011111" => valeur <= X"0D0C";
		when "0010100000" => valeur <= X"0D1F";
		when "0010100001" => valeur <= X"0D33";
		when "0010100010" => valeur <= X"0D46";
		when "0010100011" => valeur <= X"0D59";
		when "0010100100" => valeur <= X"0D6C";
		when "0010100101" => valeur <= X"0D7F";
		when "0010100110" => valeur <= X"0D92";
		when "0010100111" => valeur <= X"0DA5";
		when "0010101000" => valeur <= X"0DB8";
		when "0010101001" => valeur <= X"0DCB";
		when "0010101010" => valeur <= X"0DDE";
		when "0010101011" => valeur <= X"0DF1";
		when "0010101100" => valeur <= X"0E04";
		when "0010101101" => valeur <= X"0E17";
		when "0010101110" => valeur <= X"0E2A";
		when "0010101111" => valeur <= X"0E3D";
		when "0010110000" => valeur <= X"0E50";
		when "0010110001" => valeur <= X"0E62";
		when "0010110010" => valeur <= X"0E75";
		when "0010110011" => valeur <= X"0E88";
		when "0010110100" => valeur <= X"0E9A";
		when "0010110101" => valeur <= X"0EAD";
		when "0010110110" => valeur <= X"0EBF";
		when "0010110111" => valeur <= X"0ED2";
		when "0010111000" => valeur <= X"0EE4";
		when "0010111001" => valeur <= X"0EF7";
		when "0010111010" => valeur <= X"0F09";
		when "0010111011" => valeur <= X"0F1C";
		when "0010111100" => valeur <= X"0F2E";
		when "0010111101" => valeur <= X"0F40";
		when "0010111110" => valeur <= X"0F53";
		when "0010111111" => valeur <= X"0F65";
		when "0011000000" => valeur <= X"0F77";
		when "0011000001" => valeur <= X"0F89";
		when "0011000010" => valeur <= X"0F9B";
		when "0011000011" => valeur <= X"0FAD";
		when "0011000100" => valeur <= X"0FBF";
		when "0011000101" => valeur <= X"0FD1";
		when "0011000110" => valeur <= X"0FE3";
		when "0011000111" => valeur <= X"0FF5";
		when "0011001000" => valeur <= X"1007";
		when "0011001001" => valeur <= X"1019";
		when "0011001010" => valeur <= X"102B";
		when "0011001011" => valeur <= X"103D";
		when "0011001100" => valeur <= X"104E";
		when "0011001101" => valeur <= X"1060";
		when "0011001110" => valeur <= X"1072";
		when "0011001111" => valeur <= X"1083";
		when "0011010000" => valeur <= X"1095";
		when "0011010001" => valeur <= X"10A6";
		when "0011010010" => valeur <= X"10B8";
		when "0011010011" => valeur <= X"10C9";
		when "0011010100" => valeur <= X"10DB";
		when "0011010101" => valeur <= X"10EC";
		when "0011010110" => valeur <= X"10FE";
		when "0011010111" => valeur <= X"110F";
		when "0011011000" => valeur <= X"1120";
		when "0011011001" => valeur <= X"1131";
		when "0011011010" => valeur <= X"1142";
		when "0011011011" => valeur <= X"1154";
		when "0011011100" => valeur <= X"1165";
		when "0011011101" => valeur <= X"1176";
		when "0011011110" => valeur <= X"1187";
		when "0011011111" => valeur <= X"1198";
		when "0011100000" => valeur <= X"11A9";
		when "0011100001" => valeur <= X"11BA";
		when "0011100010" => valeur <= X"11CA";
		when "0011100011" => valeur <= X"11DB";
		when "0011100100" => valeur <= X"11EC";
		when "0011100101" => valeur <= X"11FD";
		when "0011100110" => valeur <= X"120D";
		when "0011100111" => valeur <= X"121E";
		when "0011101000" => valeur <= X"122E";
		when "0011101001" => valeur <= X"123F";
		when "0011101010" => valeur <= X"124F";
		when "0011101011" => valeur <= X"1260";
		when "0011101100" => valeur <= X"1270";
		when "0011101101" => valeur <= X"1281";
		when "0011101110" => valeur <= X"1291";
		when "0011101111" => valeur <= X"12A1";
		when "0011110000" => valeur <= X"12B1";
		when "0011110001" => valeur <= X"12C2";
		when "0011110010" => valeur <= X"12D2";
		when "0011110011" => valeur <= X"12E2";
		when "0011110100" => valeur <= X"12F2";
		when "0011110101" => valeur <= X"1302";
		when "0011110110" => valeur <= X"1312";
		when "0011110111" => valeur <= X"1322";
		when "0011111000" => valeur <= X"1332";
		when "0011111001" => valeur <= X"1341";
		when "0011111010" => valeur <= X"1351";
		when "0011111011" => valeur <= X"1361";
		when "0011111100" => valeur <= X"1370";
		when "0011111101" => valeur <= X"1380";
		when "0011111110" => valeur <= X"1390";
		when "0011111111" => valeur <= X"139F";
		when "0100000000" => valeur <= X"13AF";
		when "0100000001" => valeur <= X"13BE";
		when "0100000010" => valeur <= X"13CD";
		when "0100000011" => valeur <= X"13DD";
		when "0100000100" => valeur <= X"13EC";
		when "0100000101" => valeur <= X"13FB";
		when "0100000110" => valeur <= X"140B";
		when "0100000111" => valeur <= X"141A";
		when "0100001000" => valeur <= X"1429";
		when "0100001001" => valeur <= X"1438";
		when "0100001010" => valeur <= X"1447";
		when "0100001011" => valeur <= X"1456";
		when "0100001100" => valeur <= X"1465";
		when "0100001101" => valeur <= X"1473";
		when "0100001110" => valeur <= X"1482";
		when "0100001111" => valeur <= X"1491";
		when "0100010000" => valeur <= X"14A0";
		when "0100010001" => valeur <= X"14AE";
		when "0100010010" => valeur <= X"14BD";
		when "0100010011" => valeur <= X"14CC";
		when "0100010100" => valeur <= X"14DA";
		when "0100010101" => valeur <= X"14E9";
		when "0100010110" => valeur <= X"14F7";
		when "0100010111" => valeur <= X"1505";
		when "0100011000" => valeur <= X"1514";
		when "0100011001" => valeur <= X"1522";
		when "0100011010" => valeur <= X"1530";
		when "0100011011" => valeur <= X"153E";
		when "0100011100" => valeur <= X"154C";
		when "0100011101" => valeur <= X"155A";
		when "0100011110" => valeur <= X"1568";
		when "0100011111" => valeur <= X"1576";
		when "0100100000" => valeur <= X"1584";
		when "0100100001" => valeur <= X"1592";
		when "0100100010" => valeur <= X"15A0";
		when "0100100011" => valeur <= X"15AD";
		when "0100100100" => valeur <= X"15BB";
		when "0100100101" => valeur <= X"15C9";
		when "0100100110" => valeur <= X"15D6";
		when "0100100111" => valeur <= X"15E4";
		when "0100101000" => valeur <= X"15F1";
		when "0100101001" => valeur <= X"15FF";
		when "0100101010" => valeur <= X"160C";
		when "0100101011" => valeur <= X"1619";
		when "0100101100" => valeur <= X"1627";
		when "0100101101" => valeur <= X"1634";
		when "0100101110" => valeur <= X"1641";
		when "0100101111" => valeur <= X"164E";
		when "0100110000" => valeur <= X"165B";
		when "0100110001" => valeur <= X"1668";
		when "0100110010" => valeur <= X"1675";
		when "0100110011" => valeur <= X"1682";
		when "0100110100" => valeur <= X"168F";
		when "0100110101" => valeur <= X"169C";
		when "0100110110" => valeur <= X"16A8";
		when "0100110111" => valeur <= X"16B5";
		when "0100111000" => valeur <= X"16C2";
		when "0100111001" => valeur <= X"16CE";
		when "0100111010" => valeur <= X"16DB";
		when "0100111011" => valeur <= X"16E7";
		when "0100111100" => valeur <= X"16F3";
		when "0100111101" => valeur <= X"1700";
		when "0100111110" => valeur <= X"170C";
		when "0100111111" => valeur <= X"1718";
		when "0101000000" => valeur <= X"1724";
		when "0101000001" => valeur <= X"1731";
		when "0101000010" => valeur <= X"173D";
		when "0101000011" => valeur <= X"1749";
		when "0101000100" => valeur <= X"1755";
		when "0101000101" => valeur <= X"1760";
		when "0101000110" => valeur <= X"176C";
		when "0101000111" => valeur <= X"1778";
		when "0101001000" => valeur <= X"1784";
		when "0101001001" => valeur <= X"178F";
		when "0101001010" => valeur <= X"179B";
		when "0101001011" => valeur <= X"17A7";
		when "0101001100" => valeur <= X"17B2";
		when "0101001101" => valeur <= X"17BD";
		when "0101001110" => valeur <= X"17C9";
		when "0101001111" => valeur <= X"17D4";
		when "0101010000" => valeur <= X"17DF";
		when "0101010001" => valeur <= X"17EB";
		when "0101010010" => valeur <= X"17F6";
		when "0101010011" => valeur <= X"1801";
		when "0101010100" => valeur <= X"180C";
		when "0101010101" => valeur <= X"1817";
		when "0101010110" => valeur <= X"1822";
		when "0101010111" => valeur <= X"182D";
		when "0101011000" => valeur <= X"1837";
		when "0101011001" => valeur <= X"1842";
		when "0101011010" => valeur <= X"184D";
		when "0101011011" => valeur <= X"1857";
		when "0101011100" => valeur <= X"1862";
		when "0101011101" => valeur <= X"186D";
		when "0101011110" => valeur <= X"1877";
		when "0101011111" => valeur <= X"1881";
		when "0101100000" => valeur <= X"188C";
		when "0101100001" => valeur <= X"1896";
		when "0101100010" => valeur <= X"18A0";
		when "0101100011" => valeur <= X"18AA";
		when "0101100100" => valeur <= X"18B4";
		when "0101100101" => valeur <= X"18BE";
		when "0101100110" => valeur <= X"18C8";
		when "0101100111" => valeur <= X"18D2";
		when "0101101000" => valeur <= X"18DC";
		when "0101101001" => valeur <= X"18E6";
		when "0101101010" => valeur <= X"18F0";
		when "0101101011" => valeur <= X"18F9";
		when "0101101100" => valeur <= X"1903";
		when "0101101101" => valeur <= X"190D";
		when "0101101110" => valeur <= X"1916";
		when "0101101111" => valeur <= X"191F";
		when "0101110000" => valeur <= X"1929";
		when "0101110001" => valeur <= X"1932";
		when "0101110010" => valeur <= X"193B";
		when "0101110011" => valeur <= X"1945";
		when "0101110100" => valeur <= X"194E";
		when "0101110101" => valeur <= X"1957";
		when "0101110110" => valeur <= X"1960";
		when "0101110111" => valeur <= X"1969";
		when "0101111000" => valeur <= X"1972";
		when "0101111001" => valeur <= X"197A";
		when "0101111010" => valeur <= X"1983";
		when "0101111011" => valeur <= X"198C";
		when "0101111100" => valeur <= X"1994";
		when "0101111101" => valeur <= X"199D";
		when "0101111110" => valeur <= X"19A6";
		when "0101111111" => valeur <= X"19AE";
		when "0110000000" => valeur <= X"19B6";
		when "0110000001" => valeur <= X"19BF";
		when "0110000010" => valeur <= X"19C7";
		when "0110000011" => valeur <= X"19CF";
		when "0110000100" => valeur <= X"19D7";
		when "0110000101" => valeur <= X"19DF";
		when "0110000110" => valeur <= X"19E7";
		when "0110000111" => valeur <= X"19EF";
		when "0110001000" => valeur <= X"19F7";
		when "0110001001" => valeur <= X"19FF";
		when "0110001010" => valeur <= X"1A07";
		when "0110001011" => valeur <= X"1A0F";
		when "0110001100" => valeur <= X"1A16";
		when "0110001101" => valeur <= X"1A1E";
		when "0110001110" => valeur <= X"1A25";
		when "0110001111" => valeur <= X"1A2D";
		when "0110010000" => valeur <= X"1A34";
		when "0110010001" => valeur <= X"1A3B";
		when "0110010010" => valeur <= X"1A43";
		when "0110010011" => valeur <= X"1A4A";
		when "0110010100" => valeur <= X"1A51";
		when "0110010101" => valeur <= X"1A58";
		when "0110010110" => valeur <= X"1A5F";
		when "0110010111" => valeur <= X"1A66";
		when "0110011000" => valeur <= X"1A6D";
		when "0110011001" => valeur <= X"1A74";
		when "0110011010" => valeur <= X"1A7A";
		when "0110011011" => valeur <= X"1A81";
		when "0110011100" => valeur <= X"1A88";
		when "0110011101" => valeur <= X"1A8E";
		when "0110011110" => valeur <= X"1A95";
		when "0110011111" => valeur <= X"1A9B";
		when "0110100000" => valeur <= X"1AA2";
		when "0110100001" => valeur <= X"1AA8";
		when "0110100010" => valeur <= X"1AAE";
		when "0110100011" => valeur <= X"1AB4";
		when "0110100100" => valeur <= X"1ABA";
		when "0110100101" => valeur <= X"1AC0";
		when "0110100110" => valeur <= X"1AC6";
		when "0110100111" => valeur <= X"1ACC";
		when "0110101000" => valeur <= X"1AD2";
		when "0110101001" => valeur <= X"1AD8";
		when "0110101010" => valeur <= X"1ADE";
		when "0110101011" => valeur <= X"1AE3";
		when "0110101100" => valeur <= X"1AE9";
		when "0110101101" => valeur <= X"1AEE";
		when "0110101110" => valeur <= X"1AF4";
		when "0110101111" => valeur <= X"1AF9";
		when "0110110000" => valeur <= X"1AFF";
		when "0110110001" => valeur <= X"1B04";
		when "0110110010" => valeur <= X"1B09";
		when "0110110011" => valeur <= X"1B0E";
		when "0110110100" => valeur <= X"1B13";
		when "0110110101" => valeur <= X"1B18";
		when "0110110110" => valeur <= X"1B1D";
		when "0110110111" => valeur <= X"1B22";
		when "0110111000" => valeur <= X"1B27";
		when "0110111001" => valeur <= X"1B2C";
		when "0110111010" => valeur <= X"1B30";
		when "0110111011" => valeur <= X"1B35";
		when "0110111100" => valeur <= X"1B3A";
		when "0110111101" => valeur <= X"1B3E";
		when "0110111110" => valeur <= X"1B42";
		when "0110111111" => valeur <= X"1B47";
		when "0111000000" => valeur <= X"1B4B";
		when "0111000001" => valeur <= X"1B4F";
		when "0111000010" => valeur <= X"1B53";
		when "0111000011" => valeur <= X"1B58";
		when "0111000100" => valeur <= X"1B5C";
		when "0111000101" => valeur <= X"1B5F";
		when "0111000110" => valeur <= X"1B63";
		when "0111000111" => valeur <= X"1B67";
		when "0111001000" => valeur <= X"1B6B";
		when "0111001001" => valeur <= X"1B6F";
		when "0111001010" => valeur <= X"1B72";
		when "0111001011" => valeur <= X"1B76";
		when "0111001100" => valeur <= X"1B79";
		when "0111001101" => valeur <= X"1B7D";
		when "0111001110" => valeur <= X"1B80";
		when "0111001111" => valeur <= X"1B83";
		when "0111010000" => valeur <= X"1B87";
		when "0111010001" => valeur <= X"1B8A";
		when "0111010010" => valeur <= X"1B8D";
		when "0111010011" => valeur <= X"1B90";
		when "0111010100" => valeur <= X"1B93";
		when "0111010101" => valeur <= X"1B96";
		when "0111010110" => valeur <= X"1B99";
		when "0111010111" => valeur <= X"1B9B";
		when "0111011000" => valeur <= X"1B9E";
		when "0111011001" => valeur <= X"1BA1";
		when "0111011010" => valeur <= X"1BA3";
		when "0111011011" => valeur <= X"1BA6";
		when "0111011100" => valeur <= X"1BA8";
		when "0111011101" => valeur <= X"1BAB";
		when "0111011110" => valeur <= X"1BAD";
		when "0111011111" => valeur <= X"1BAF";
		when "0111100000" => valeur <= X"1BB1";
		when "0111100001" => valeur <= X"1BB3";
		when "0111100010" => valeur <= X"1BB5";
		when "0111100011" => valeur <= X"1BB7";
		when "0111100100" => valeur <= X"1BB9";
		when "0111100101" => valeur <= X"1BBB";
		when "0111100110" => valeur <= X"1BBD";
		when "0111100111" => valeur <= X"1BBE";
		when "0111101000" => valeur <= X"1BC0";
		when "0111101001" => valeur <= X"1BC2";
		when "0111101010" => valeur <= X"1BC3";
		when "0111101011" => valeur <= X"1BC5";
		when "0111101100" => valeur <= X"1BC6";
		when "0111101101" => valeur <= X"1BC7";
		when "0111101110" => valeur <= X"1BC8";
		when "0111101111" => valeur <= X"1BCA";
		when "0111110000" => valeur <= X"1BCB";
		when "0111110001" => valeur <= X"1BCC";
		when "0111110010" => valeur <= X"1BCD";
		when "0111110011" => valeur <= X"1BCE";
		when "0111110100" => valeur <= X"1BCE";
		when "0111110101" => valeur <= X"1BCF";
		when "0111110110" => valeur <= X"1BD0";
		when "0111110111" => valeur <= X"1BD0";
		when "0111111000" => valeur <= X"1BD1";
		when "0111111001" => valeur <= X"1BD1";
		when "0111111010" => valeur <= X"1BD2";
		when "0111111011" => valeur <= X"1BD2";
		when "0111111100" => valeur <= X"1BD3";
		when "0111111101" => valeur <= X"1BD3";
		when "0111111110" => valeur <= X"1BD3";
		when "0111111111" => valeur <= X"1BD3";
		when "1000000000" => valeur <= X"1BD3";
		when "1000000001" => valeur <= X"1BD3";
		when "1000000010" => valeur <= X"1BD3";
		when "1000000011" => valeur <= X"1BD3";
		when "1000000100" => valeur <= X"1BD2";
		when "1000000101" => valeur <= X"1BD2";
		when "1000000110" => valeur <= X"1BD2";
		when "1000000111" => valeur <= X"1BD1";
		when "1000001000" => valeur <= X"1BD1";
		when "1000001001" => valeur <= X"1BD0";
		when "1000001010" => valeur <= X"1BCF";
		when "1000001011" => valeur <= X"1BCF";
		when "1000001100" => valeur <= X"1BCE";
		when "1000001101" => valeur <= X"1BCD";
		when "1000001110" => valeur <= X"1BCC";
		when "1000001111" => valeur <= X"1BCB";
		when "1000010000" => valeur <= X"1BCA";
		when "1000010001" => valeur <= X"1BC9";
		when "1000010010" => valeur <= X"1BC8";
		when "1000010011" => valeur <= X"1BC7";
		when "1000010100" => valeur <= X"1BC5";
		when "1000010101" => valeur <= X"1BC4";
		when "1000010110" => valeur <= X"1BC2";
		when "1000010111" => valeur <= X"1BC1";
		when "1000011000" => valeur <= X"1BBF";
		when "1000011001" => valeur <= X"1BBE";
		when "1000011010" => valeur <= X"1BBC";
		when "1000011011" => valeur <= X"1BBA";
		when "1000011100" => valeur <= X"1BB8";
		when "1000011101" => valeur <= X"1BB6";
		when "1000011110" => valeur <= X"1BB4";
		when "1000011111" => valeur <= X"1BB2";
		when "1000100000" => valeur <= X"1BB0";
		when "1000100001" => valeur <= X"1BAE";
		when "1000100010" => valeur <= X"1BAC";
		when "1000100011" => valeur <= X"1BA9";
		when "1000100100" => valeur <= X"1BA7";
		when "1000100101" => valeur <= X"1BA4";
		when "1000100110" => valeur <= X"1BA2";
		when "1000100111" => valeur <= X"1B9F";
		when "1000101000" => valeur <= X"1B9D";
		when "1000101001" => valeur <= X"1B9A";
		when "1000101010" => valeur <= X"1B97";
		when "1000101011" => valeur <= X"1B94";
		when "1000101100" => valeur <= X"1B91";
		when "1000101101" => valeur <= X"1B8E";
		when "1000101110" => valeur <= X"1B8B";
		when "1000101111" => valeur <= X"1B88";
		when "1000110000" => valeur <= X"1B85";
		when "1000110001" => valeur <= X"1B82";
		when "1000110010" => valeur <= X"1B7E";
		when "1000110011" => valeur <= X"1B7B";
		when "1000110100" => valeur <= X"1B78";
		when "1000110101" => valeur <= X"1B74";
		when "1000110110" => valeur <= X"1B70";
		when "1000110111" => valeur <= X"1B6D";
		when "1000111000" => valeur <= X"1B69";
		when "1000111001" => valeur <= X"1B65";
		when "1000111010" => valeur <= X"1B61";
		when "1000111011" => valeur <= X"1B5E";
		when "1000111100" => valeur <= X"1B5A";
		when "1000111101" => valeur <= X"1B55";
		when "1000111110" => valeur <= X"1B51";
		when "1000111111" => valeur <= X"1B4D";
		when "1001000000" => valeur <= X"1B49";
		when "1001000001" => valeur <= X"1B45";
		when "1001000010" => valeur <= X"1B40";
		when "1001000011" => valeur <= X"1B3C";
		when "1001000100" => valeur <= X"1B37";
		when "1001000101" => valeur <= X"1B33";
		when "1001000110" => valeur <= X"1B2E";
		when "1001000111" => valeur <= X"1B29";
		when "1001001000" => valeur <= X"1B25";
		when "1001001001" => valeur <= X"1B20";
		when "1001001010" => valeur <= X"1B1B";
		when "1001001011" => valeur <= X"1B16";
		when "1001001100" => valeur <= X"1B11";
		when "1001001101" => valeur <= X"1B0C";
		when "1001001110" => valeur <= X"1B07";
		when "1001001111" => valeur <= X"1B01";
		when "1001010000" => valeur <= X"1AFC";
		when "1001010001" => valeur <= X"1AF7";
		when "1001010010" => valeur <= X"1AF1";
		when "1001010011" => valeur <= X"1AEC";
		when "1001010100" => valeur <= X"1AE6";
		when "1001010101" => valeur <= X"1AE1";
		when "1001010110" => valeur <= X"1ADB";
		when "1001010111" => valeur <= X"1AD5";
		when "1001011000" => valeur <= X"1ACF";
		when "1001011001" => valeur <= X"1AC9";
		when "1001011010" => valeur <= X"1AC3";
		when "1001011011" => valeur <= X"1ABD";
		when "1001011100" => valeur <= X"1AB7";
		when "1001011101" => valeur <= X"1AB1";
		when "1001011110" => valeur <= X"1AAB";
		when "1001011111" => valeur <= X"1AA5";
		when "1001100000" => valeur <= X"1A9E";
		when "1001100001" => valeur <= X"1A98";
		when "1001100010" => valeur <= X"1A92";
		when "1001100011" => valeur <= X"1A8B";
		when "1001100100" => valeur <= X"1A84";
		when "1001100101" => valeur <= X"1A7E";
		when "1001100110" => valeur <= X"1A77";
		when "1001100111" => valeur <= X"1A70";
		when "1001101000" => valeur <= X"1A69";
		when "1001101001" => valeur <= X"1A63";
		when "1001101010" => valeur <= X"1A5C";
		when "1001101011" => valeur <= X"1A55";
		when "1001101100" => valeur <= X"1A4D";
		when "1001101101" => valeur <= X"1A46";
		when "1001101110" => valeur <= X"1A3F";
		when "1001101111" => valeur <= X"1A38";
		when "1001110000" => valeur <= X"1A30";
		when "1001110001" => valeur <= X"1A29";
		when "1001110010" => valeur <= X"1A21";
		when "1001110011" => valeur <= X"1A1A";
		when "1001110100" => valeur <= X"1A12";
		when "1001110101" => valeur <= X"1A0B";
		when "1001110110" => valeur <= X"1A03";
		when "1001110111" => valeur <= X"19FB";
		when "1001111000" => valeur <= X"19F3";
		when "1001111001" => valeur <= X"19EB";
		when "1001111010" => valeur <= X"19E3";
		when "1001111011" => valeur <= X"19DB";
		when "1001111100" => valeur <= X"19D3";
		when "1001111101" => valeur <= X"19CB";
		when "1001111110" => valeur <= X"19C3";
		when "1001111111" => valeur <= X"19BB";
		when "1010000000" => valeur <= X"19B2";
		when "1010000001" => valeur <= X"19AA";
		when "1010000010" => valeur <= X"19A1";
		when "1010000011" => valeur <= X"1999";
		when "1010000100" => valeur <= X"1990";
		when "1010000101" => valeur <= X"1987";
		when "1010000110" => valeur <= X"197F";
		when "1010000111" => valeur <= X"1976";
		when "1010001000" => valeur <= X"196D";
		when "1010001001" => valeur <= X"1964";
		when "1010001010" => valeur <= X"195B";
		when "1010001011" => valeur <= X"1952";
		when "1010001100" => valeur <= X"1949";
		when "1010001101" => valeur <= X"1940";
		when "1010001110" => valeur <= X"1937";
		when "1010001111" => valeur <= X"192D";
		when "1010010000" => valeur <= X"1924";
		when "1010010001" => valeur <= X"191B";
		when "1010010010" => valeur <= X"1911";
		when "1010010011" => valeur <= X"1908";
		when "1010010100" => valeur <= X"18FE";
		when "1010010101" => valeur <= X"18F5";
		when "1010010110" => valeur <= X"18EB";
		when "1010010111" => valeur <= X"18E1";
		when "1010011000" => valeur <= X"18D7";
		when "1010011001" => valeur <= X"18CD";
		when "1010011010" => valeur <= X"18C3";
		when "1010011011" => valeur <= X"18B9";
		when "1010011100" => valeur <= X"18AF";
		when "1010011101" => valeur <= X"18A5";
		when "1010011110" => valeur <= X"189B";
		when "1010011111" => valeur <= X"1891";
		when "1010100000" => valeur <= X"1887";
		when "1010100001" => valeur <= X"187C";
		when "1010100010" => valeur <= X"1872";
		when "1010100011" => valeur <= X"1867";
		when "1010100100" => valeur <= X"185D";
		when "1010100101" => valeur <= X"1852";
		when "1010100110" => valeur <= X"1848";
		when "1010100111" => valeur <= X"183D";
		when "1010101000" => valeur <= X"1832";
		when "1010101001" => valeur <= X"1827";
		when "1010101010" => valeur <= X"181C";
		when "1010101011" => valeur <= X"1811";
		when "1010101100" => valeur <= X"1806";
		when "1010101101" => valeur <= X"17FB";
		when "1010101110" => valeur <= X"17F0";
		when "1010101111" => valeur <= X"17E5";
		when "1010110000" => valeur <= X"17DA";
		when "1010110001" => valeur <= X"17CF";
		when "1010110010" => valeur <= X"17C3";
		when "1010110011" => valeur <= X"17B8";
		when "1010110100" => valeur <= X"17AC";
		when "1010110101" => valeur <= X"17A1";
		when "1010110110" => valeur <= X"1795";
		when "1010110111" => valeur <= X"178A";
		when "1010111000" => valeur <= X"177E";
		when "1010111001" => valeur <= X"1772";
		when "1010111010" => valeur <= X"1766";
		when "1010111011" => valeur <= X"175B";
		when "1010111100" => valeur <= X"174F";
		when "1010111101" => valeur <= X"1743";
		when "1010111110" => valeur <= X"1737";
		when "1010111111" => valeur <= X"172B";
		when "1011000000" => valeur <= X"171E";
		when "1011000001" => valeur <= X"1712";
		when "1011000010" => valeur <= X"1706";
		when "1011000011" => valeur <= X"16FA";
		when "1011000100" => valeur <= X"16ED";
		when "1011000101" => valeur <= X"16E1";
		when "1011000110" => valeur <= X"16D4";
		when "1011000111" => valeur <= X"16C8";
		when "1011001000" => valeur <= X"16BB";
		when "1011001001" => valeur <= X"16AF";
		when "1011001010" => valeur <= X"16A2";
		when "1011001011" => valeur <= X"1695";
		when "1011001100" => valeur <= X"1688";
		when "1011001101" => valeur <= X"167C";
		when "1011001110" => valeur <= X"166F";
		when "1011001111" => valeur <= X"1662";
		when "1011010000" => valeur <= X"1655";
		when "1011010001" => valeur <= X"1648";
		when "1011010010" => valeur <= X"163A";
		when "1011010011" => valeur <= X"162D";
		when "1011010100" => valeur <= X"1620";
		when "1011010101" => valeur <= X"1613";
		when "1011010110" => valeur <= X"1605";
		when "1011010111" => valeur <= X"15F8";
		when "1011011000" => valeur <= X"15EB";
		when "1011011001" => valeur <= X"15DD";
		when "1011011010" => valeur <= X"15D0";
		when "1011011011" => valeur <= X"15C2";
		when "1011011100" => valeur <= X"15B4";
		when "1011011101" => valeur <= X"15A7";
		when "1011011110" => valeur <= X"1599";
		when "1011011111" => valeur <= X"158B";
		when "1011100000" => valeur <= X"157D";
		when "1011100001" => valeur <= X"156F";
		when "1011100010" => valeur <= X"1561";
		when "1011100011" => valeur <= X"1553";
		when "1011100100" => valeur <= X"1545";
		when "1011100101" => valeur <= X"1537";
		when "1011100110" => valeur <= X"1529";
		when "1011100111" => valeur <= X"151B";
		when "1011101000" => valeur <= X"150C";
		when "1011101001" => valeur <= X"14FE";
		when "1011101010" => valeur <= X"14F0";
		when "1011101011" => valeur <= X"14E1";
		when "1011101100" => valeur <= X"14D3";
		when "1011101101" => valeur <= X"14C4";
		when "1011101110" => valeur <= X"14B6";
		when "1011101111" => valeur <= X"14A7";
		when "1011110000" => valeur <= X"1498";
		when "1011110001" => valeur <= X"148A";
		when "1011110010" => valeur <= X"147B";
		when "1011110011" => valeur <= X"146C";
		when "1011110100" => valeur <= X"145D";
		when "1011110101" => valeur <= X"144E";
		when "1011110110" => valeur <= X"143F";
		when "1011110111" => valeur <= X"1430";
		when "1011111000" => valeur <= X"1421";
		when "1011111001" => valeur <= X"1412";
		when "1011111010" => valeur <= X"1403";
		when "1011111011" => valeur <= X"13F4";
		when "1011111100" => valeur <= X"13E4";
		when "1011111101" => valeur <= X"13D5";
		when "1011111110" => valeur <= X"13C6";
		when "1011111111" => valeur <= X"13B6";
		when "1100000000" => valeur <= X"13A7";
		when "1100000001" => valeur <= X"1397";
		when "1100000010" => valeur <= X"1388";
		when "1100000011" => valeur <= X"1378";
		when "1100000100" => valeur <= X"1369";
		when "1100000101" => valeur <= X"1359";
		when "1100000110" => valeur <= X"1349";
		when "1100000111" => valeur <= X"1339";
		when "1100001000" => valeur <= X"132A";
		when "1100001001" => valeur <= X"131A";
		when "1100001010" => valeur <= X"130A";
		when "1100001011" => valeur <= X"12FA";
		when "1100001100" => valeur <= X"12EA";
		when "1100001101" => valeur <= X"12DA";
		when "1100001110" => valeur <= X"12CA";
		when "1100001111" => valeur <= X"12BA";
		when "1100010000" => valeur <= X"12A9";
		when "1100010001" => valeur <= X"1299";
		when "1100010010" => valeur <= X"1289";
		when "1100010011" => valeur <= X"1278";
		when "1100010100" => valeur <= X"1268";
		when "1100010101" => valeur <= X"1258";
		when "1100010110" => valeur <= X"1247";
		when "1100010111" => valeur <= X"1237";
		when "1100011000" => valeur <= X"1226";
		when "1100011001" => valeur <= X"1216";
		when "1100011010" => valeur <= X"1205";
		when "1100011011" => valeur <= X"11F4";
		when "1100011100" => valeur <= X"11E4";
		when "1100011101" => valeur <= X"11D3";
		when "1100011110" => valeur <= X"11C2";
		when "1100011111" => valeur <= X"11B1";
		when "1100100000" => valeur <= X"11A0";
		when "1100100001" => valeur <= X"118F";
		when "1100100010" => valeur <= X"117E";
		when "1100100011" => valeur <= X"116D";
		when "1100100100" => valeur <= X"115C";
		when "1100100101" => valeur <= X"114B";
		when "1100100110" => valeur <= X"113A";
		when "1100100111" => valeur <= X"1129";
		when "1100101000" => valeur <= X"1117";
		when "1100101001" => valeur <= X"1106";
		when "1100101010" => valeur <= X"10F5";
		when "1100101011" => valeur <= X"10E4";
		when "1100101100" => valeur <= X"10D2";
		when "1100101101" => valeur <= X"10C1";
		when "1100101110" => valeur <= X"10AF";
		when "1100101111" => valeur <= X"109E";
		when "1100110000" => valeur <= X"108C";
		when "1100110001" => valeur <= X"107B";
		when "1100110010" => valeur <= X"1069";
		when "1100110011" => valeur <= X"1057";
		when "1100110100" => valeur <= X"1046";
		when "1100110101" => valeur <= X"1034";
		when "1100110110" => valeur <= X"1022";
		when "1100110111" => valeur <= X"1010";
		when "1100111000" => valeur <= X"0FFE";
		when "1100111001" => valeur <= X"0FEC";
		when "1100111010" => valeur <= X"0FDA";
		when "1100111011" => valeur <= X"0FC8";
		when "1100111100" => valeur <= X"0FB6";
		when "1100111101" => valeur <= X"0FA4";
		when "1100111110" => valeur <= X"0F92";
		when "1100111111" => valeur <= X"0F80";
		when "1101000000" => valeur <= X"0F6E";
		when "1101000001" => valeur <= X"0F5C";
		when "1101000010" => valeur <= X"0F49";
		when "1101000011" => valeur <= X"0F37";
		when "1101000100" => valeur <= X"0F25";
		when "1101000101" => valeur <= X"0F13";
		when "1101000110" => valeur <= X"0F00";
		when "1101000111" => valeur <= X"0EEE";
		when "1101001000" => valeur <= X"0EDB";
		when "1101001001" => valeur <= X"0EC9";
		when "1101001010" => valeur <= X"0EB6";
		when "1101001011" => valeur <= X"0EA4";
		when "1101001100" => valeur <= X"0E91";
		when "1101001101" => valeur <= X"0E7E";
		when "1101001110" => valeur <= X"0E6C";
		when "1101001111" => valeur <= X"0E59";
		when "1101010000" => valeur <= X"0E46";
		when "1101010001" => valeur <= X"0E33";
		when "1101010010" => valeur <= X"0E21";
		when "1101010011" => valeur <= X"0E0E";
		when "1101010100" => valeur <= X"0DFB";
		when "1101010101" => valeur <= X"0DE8";
		when "1101010110" => valeur <= X"0DD5";
		when "1101010111" => valeur <= X"0DC2";
		when "1101011000" => valeur <= X"0DAF";
		when "1101011001" => valeur <= X"0D9C";
		when "1101011010" => valeur <= X"0D89";
		when "1101011011" => valeur <= X"0D76";
		when "1101011100" => valeur <= X"0D63";
		when "1101011101" => valeur <= X"0D4F";
		when "1101011110" => valeur <= X"0D3C";
		when "1101011111" => valeur <= X"0D29";
		when "1101100000" => valeur <= X"0D16";
		when "1101100001" => valeur <= X"0D02";
		when "1101100010" => valeur <= X"0CEF";
		when "1101100011" => valeur <= X"0CDC";
		when "1101100100" => valeur <= X"0CC8";
		when "1101100101" => valeur <= X"0CB5";
		when "1101100110" => valeur <= X"0CA1";
		when "1101100111" => valeur <= X"0C8E";
		when "1101101000" => valeur <= X"0C7A";
		when "1101101001" => valeur <= X"0C67";
		when "1101101010" => valeur <= X"0C53";
		when "1101101011" => valeur <= X"0C40";
		when "1101101100" => valeur <= X"0C2C";
		when "1101101101" => valeur <= X"0C18";
		when "1101101110" => valeur <= X"0C04";
		when "1101101111" => valeur <= X"0BF1";
		when "1101110000" => valeur <= X"0BDD";
		when "1101110001" => valeur <= X"0BC9";
		when "1101110010" => valeur <= X"0BB5";
		when "1101110011" => valeur <= X"0BA2";
		when "1101110100" => valeur <= X"0B8E";
		when "1101110101" => valeur <= X"0B7A";
		when "1101110110" => valeur <= X"0B66";
		when "1101110111" => valeur <= X"0B52";
		when "1101111000" => valeur <= X"0B3E";
		when "1101111001" => valeur <= X"0B2A";
		when "1101111010" => valeur <= X"0B16";
		when "1101111011" => valeur <= X"0B02";
		when "1101111100" => valeur <= X"0AEE";
		when "1101111101" => valeur <= X"0ADA";
		when "1101111110" => valeur <= X"0AC5";
		when "1101111111" => valeur <= X"0AB1";
		when "1110000000" => valeur <= X"0A9D";
		when "1110000001" => valeur <= X"0A89";
		when "1110000010" => valeur <= X"0A75";
		when "1110000011" => valeur <= X"0A60";
		when "1110000100" => valeur <= X"0A4C";
		when "1110000101" => valeur <= X"0A38";
		when "1110000110" => valeur <= X"0A23";
		when "1110000111" => valeur <= X"0A0F";
		when "1110001000" => valeur <= X"09FB";
		when "1110001001" => valeur <= X"09E6";
		when "1110001010" => valeur <= X"09D2";
		when "1110001011" => valeur <= X"09BD";
		when "1110001100" => valeur <= X"09A9";
		when "1110001101" => valeur <= X"0994";
		when "1110001110" => valeur <= X"0980";
		when "1110001111" => valeur <= X"096B";
		when "1110010000" => valeur <= X"0956";
		when "1110010001" => valeur <= X"0942";
		when "1110010010" => valeur <= X"092D";
		when "1110010011" => valeur <= X"0919";
		when "1110010100" => valeur <= X"0904";
		when "1110010101" => valeur <= X"08EF";
		when "1110010110" => valeur <= X"08DB";
		when "1110010111" => valeur <= X"08C6";
		when "1110011000" => valeur <= X"08B1";
		when "1110011001" => valeur <= X"089C";
		when "1110011010" => valeur <= X"0887";
		when "1110011011" => valeur <= X"0873";
		when "1110011100" => valeur <= X"085E";
		when "1110011101" => valeur <= X"0849";
		when "1110011110" => valeur <= X"0834";
		when "1110011111" => valeur <= X"081F";
		when "1110100000" => valeur <= X"080A";
		when "1110100001" => valeur <= X"07F5";
		when "1110100010" => valeur <= X"07E0";
		when "1110100011" => valeur <= X"07CB";
		when "1110100100" => valeur <= X"07B6";
		when "1110100101" => valeur <= X"07A1";
		when "1110100110" => valeur <= X"078C";
		when "1110100111" => valeur <= X"0777";
		when "1110101000" => valeur <= X"0762";
		when "1110101001" => valeur <= X"074D";
		when "1110101010" => valeur <= X"0738";
		when "1110101011" => valeur <= X"0723";
		when "1110101100" => valeur <= X"070E";
		when "1110101101" => valeur <= X"06F9";
		when "1110101110" => valeur <= X"06E3";
		when "1110101111" => valeur <= X"06CE";
		when "1110110000" => valeur <= X"06B9";
		when "1110110001" => valeur <= X"06A4";
		when "1110110010" => valeur <= X"068F";
		when "1110110011" => valeur <= X"0679";
		when "1110110100" => valeur <= X"0664";
		when "1110110101" => valeur <= X"064F";
		when "1110110110" => valeur <= X"0639";
		when "1110110111" => valeur <= X"0624";
		when "1110111000" => valeur <= X"060F";
		when "1110111001" => valeur <= X"05F9";
		when "1110111010" => valeur <= X"05E4";
		when "1110111011" => valeur <= X"05CF";
		when "1110111100" => valeur <= X"05B9";
		when "1110111101" => valeur <= X"05A4";
		when "1110111110" => valeur <= X"058E";
		when "1110111111" => valeur <= X"0579";
		when "1111000000" => valeur <= X"0564";
		when "1111000001" => valeur <= X"054E";
		when "1111000010" => valeur <= X"0539";
		when "1111000011" => valeur <= X"0523";
		when "1111000100" => valeur <= X"050E";
		when "1111000101" => valeur <= X"04F8";
		when "1111000110" => valeur <= X"04E3";
		when "1111000111" => valeur <= X"04CD";
		when "1111001000" => valeur <= X"04B8";
		when "1111001001" => valeur <= X"04A2";
		when "1111001010" => valeur <= X"048C";
		when "1111001011" => valeur <= X"0477";
		when "1111001100" => valeur <= X"0461";
		when "1111001101" => valeur <= X"044C";
		when "1111001110" => valeur <= X"0436";
		when "1111001111" => valeur <= X"0420";
		when "1111010000" => valeur <= X"040B";
		when "1111010001" => valeur <= X"03F5";
		when "1111010010" => valeur <= X"03E0";
		when "1111010011" => valeur <= X"03CA";
		when "1111010100" => valeur <= X"03B4";
		when "1111010101" => valeur <= X"039F";
		when "1111010110" => valeur <= X"0389";
		when "1111010111" => valeur <= X"0373";
		when "1111011000" => valeur <= X"035E";
		when "1111011001" => valeur <= X"0348";
		when "1111011010" => valeur <= X"0332";
		when "1111011011" => valeur <= X"031C";
		when "1111011100" => valeur <= X"0307";
		when "1111011101" => valeur <= X"02F1";
		when "1111011110" => valeur <= X"02DB";
		when "1111011111" => valeur <= X"02C5";
		when "1111100000" => valeur <= X"02B0";
		when "1111100001" => valeur <= X"029A";
		when "1111100010" => valeur <= X"0284";
		when "1111100011" => valeur <= X"026E";
		when "1111100100" => valeur <= X"0259";
		when "1111100101" => valeur <= X"0243";
		when "1111100110" => valeur <= X"022D";
		when "1111100111" => valeur <= X"0217";
		when "1111101000" => valeur <= X"0201";
		when "1111101001" => valeur <= X"01EC";
		when "1111101010" => valeur <= X"01D6";
		when "1111101011" => valeur <= X"01C0";
		when "1111101100" => valeur <= X"01AA";
		when "1111101101" => valeur <= X"0194";
		when "1111101110" => valeur <= X"017E";
		when "1111101111" => valeur <= X"0169";
		when "1111110000" => valeur <= X"0153";
		when "1111110001" => valeur <= X"013D";
		when "1111110010" => valeur <= X"0127";
		when "1111110011" => valeur <= X"0111";
		when "1111110100" => valeur <= X"00FB";
		when "1111110101" => valeur <= X"00E6";
		when "1111110110" => valeur <= X"00D0";
		when "1111110111" => valeur <= X"00BA";
		when "1111111000" => valeur <= X"00A4";
		when "1111111001" => valeur <= X"008E";
		when "1111111010" => valeur <= X"0078";
		when "1111111011" => valeur <= X"0062";
		when "1111111100" => valeur <= X"004D";
		when "1111111101" => valeur <= X"0037";
		when "1111111110" => valeur <= X"0021";
		when "1111111111" => valeur <= X"000B";

		when others => valeur <= (others => '0');
	end case;
end process;
end Behavioral;

